//===========================================================================
// Module name: led_test.v
// 鏡扴: 藩路1鏃甡棒萸鏢羲楷啣奻腔LED0~LED4
//===========================================================================
`timescale 1ns / 1ps

module led_test (
                  clk,           // 羲楷啣奻怀�輮敔�: 50Mhz
                  rst_n,         // 羲楷啣奻怀�賳棒趕智�
                  led            // 怀堤LED腑,蚚衾諷秶羲楷啣奻侐跺LED(LED1~LED4)
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output [3:0] led;

//敵湔�鰶例�
reg [31:0] timer;                  
reg [3:0] led;


//===========================================================================
// 數杅�鷐�杅:悜遠數杅0~4鏃
//===========================================================================
  always @(posedge clk or negedge rst_n)    //潰聆奀笘腔奻汔朓睿葩弇腔狟蔥朓
    begin
      if (~rst_n)                           //葩弇陓瘍腴衄虴
          timer <= 0;                       //數杅�麶斲�
      else if (timer == 32'd199_999_999)    //羲楷啣妏蚚腔儒淥峈50MHzㄛ4鏃數杅(50M*4-1=199_999_999)
          timer <= 0;                       //數杅�鷐�善4鏃ㄛ數杅�麶斲�
      else
		    timer <= timer + 1'b1;            //數杅�鷐�1
    end

//===========================================================================
// LED腑諷秶
//===========================================================================
  always @(posedge clk or negedge rst_n)   //潰聆奀笘腔奻汔朓睿葩弇腔狟蔥朓
    begin
      if (~rst_n)                          //葩弇陓瘍腴衄虴
          led <= 4'b1111;                  //LED腑怀堤�屋疙舝畋譫觺ED腑謠           
      else if (timer == 32'd49_999_999)    //數杅�鷐�善1鏃ㄛ
          led <= 4'b1110;                  //LED1萸鏢
      else if (timer == 32'd99_999_999)    //數杅�鷐�善2鏃ㄛ
          led <= 4'b1101;                  //LED2萸鏢
      else if (timer == 32'd149_999_999)   //數杅�鷐�善3鏃ㄛ
          led <= 4'b1011;                  //LED3萸鏢                           
      else if (timer == 32'd199_999_999)   //數杅�鷐�善4鏃ㄛ
          led <= 4'b0111;                  //LED4萸鏢        
    end
    
endmodule

